----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/25/2022 02:21:11 PM
-- Design Name: 
-- Module Name: MPG - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- rol: sa elimine sunetul creat de buton
-- rol: sa genereze doar un sg puls (oricat as tine apasat butonul, el tot un puls va genera)

entity MPG is
    Port ( btn : in std_logic;
           clk : in std_logic;
           en : out std_logic);
end MPG;

architecture Behavioral of MPG is

Signal cnt:std_logic_vector(15 downto 0):=x"0000";
Signal Q1:std_logic := '0';
Signal Q2:std_logic := '0';
Signal Q3:std_logic := '0';

begin
    en <= Q2 AND (NOT Q3);
    
    process (clk)
    begin
        if clk'event and clk = '1' then
            cnt <= cnt + 1;
        end if;
    end process;
    
    process (clk)
    begin
        if clk'event and clk = '1' then
            if cnt(15 downto 0) = "1111111111111111" then
                Q1 <= btn;
            end if;
        end if;
    end process;
    
    process (clk)
    begin
        if clk'event and clk = '1' then
            Q2 <= Q1;
            Q3 <= Q2;
        end if;
    end process;

end Behavioral;
